module sha256_test(
	input wire clk,
	input wire data,
	output wire [255:0]result
);

sha256_transform s0(
		.state_in( 256'h5be0cd191f83d9ab9b05688c510e527fa54ff53a3c6ef372bb67ae856a09e667 ),
		.data_in( 512'h66656463626139383736353433323130666564636261393837363534333231306665646362613938373635343332313066656463626139383736353433323130 ),
		.state_out(result)
	);

endmodule
